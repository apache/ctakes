// CUI|TUI|Text|preferredTerm
C0201838|T059|Albumin
C0202202|T059|Protein
C0201850|T059|alkaline phosphatase|Alkaline phosphatase measurement
C0201836|T059|ALT|Alanine aminotransferase measurement
C0201899|T059|AST|Aspartate aminotransferase measurement
C0201913|T059|bilirubin|Bilirubin, total measurement
C0036808|T059|Bilirubin, Indirect
C0858048|T059|Bilirubin, Direct
C0201973|T059|Total CK
C0523584|T059|CK-MB|Creatine kinase MB measurement
C0523584|T059|CKMB|Creatine kinase MB measurement
C0023508|T060|white count|White Blood Cell Count procedure
C0201803|T059|osmolality|Osmolality Measurement
C0017564|T060|GFR|Glomerular Filtration Rate
C0588466|T059|RBC, UA|Red blood cells urine (lab test)
C0000010|T059|WBC, UA|White blood cells urine (lab test)
C0201837|T201|A/G Ratio|Albumin/Globulin ratio
C0373670|T059|Lipase|Lipase measurement
C0033707|T059|Protime|Prothrombin time assay
C0525032|T059|INR|International Normalized Ratio
C1443182|T059|Calc|Calculated (procedure)
C00337443|T059|sodium|Sodium measurement
C00202194|T059|potassium|Potassium measurement
C00003074|T201|Anion Gap
C00202230|T059|TSH|Thyroid stimulating hormone measurement
C01171408|T059|LDL/HDL|High density/low density lipoprotein ratio measurement
C00518015|T059|hemoglobin|Hemoglobin measurement
C00032181|T059|platelet count|Platelet Count measurement
C00018935|T059|hematocrit|Hematocrit procedure
C00201657|T059|CRP|C-reactive protein measurement
C01535922|T059|procalcitonin|Procalcitonin measurement
C00202115|T059|lactate|Lactic acid measurement
C00202225|T059|free T4|T4 free measurement
C00201934|T059|cardiac enzymes|Cardiac enzymes measurement
C00337438|T059|glucose|Glucose measurement
C00201802|T059|specific gravity|Specific gravity measurement
C00200635|T059|lymphocytes|Lymphocyte Count measurement
C00005845|T059|BUN|Blood urea nitrogen measurement
C00201975|T059|creatinine|Creatinine measurement
C01305866|T060|weight|Weighing patient
C01305855|T201|BMI|Body mass index

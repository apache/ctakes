1|1
// line comments can start with double-slash
2|3
# line comments can start with hash
3|5
4|5
C5|5
6|5
9|5
10|T5

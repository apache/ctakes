textPathFullText||^[\t ]*<Item naaccrId="textPathFullText">||<\/Item>
textPathFormalDx||^[\t ]*<Item naaccrId="textPathFormalDx">||<\/Item>
textPathClinicalHistory||^[\t ]*<Item naaccrId="textPathClinicalHistory">||<\/Item>
textDxProcPath||^[\t ]*<Item naaccrId="textDxProcPath">||<\/Item>
textPrimarySiteTitle||^[\t ]*<Item naaccrId="textPrimarySiteTitle">||<\/Item>
textHistologyTitle||^[\t ]*<Item naaccrId="textHistologyTitle">||<\/Item>
textStaging||^[\t ]*<Item naaccrId="textStaging">||<\/Item>
